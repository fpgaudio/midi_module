`ifndef __GLOBALS__
`define __GLOBALS__

// UVM Globals
localparam IN_FILE_NAME = "../tb/binary.txt";
localparam OUT_FILE_NAME = "../tb/midi.txt";
localparam CMP_FILE_NAME = "../tb/output.txt";

localparam CLK_PERIOD = 20;
localparam MIDI_CLK_PERIOD = 32000;

`endif
